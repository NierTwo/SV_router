       #       @??0��   E : \ l a b 0 \ t b . s v   