       �      �[uJ���   E : \ w 4 l a b \ t b . s v   