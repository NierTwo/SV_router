module moduleName;
    
endmodule