program automatic test(router_io.TB rtr_io);

    
endprogram